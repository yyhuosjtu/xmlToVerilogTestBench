`timescale 1ns/1ps
module PE_tb();
  parameter CYCLE=10;
  reg clk;
  reg rst;


  integer i;
  integer filez;
//pe38输出端口定义
  reg  [35:0]    PE38_Inport1;
  reg  [32:0]    PE38_Configure_Inport;
  wire [35:0]    PE38_Outport0;
  wire Pre_PE38_Bp0;
  wire Pre_PE38_Bp1;
  wire Pre_PE38_Bp2;
//end pe38 端口定义

//pe0输出端口定义
  reg  [32:0]    PE0_Configure_Inport;
  wire [35:0]    PE0_Outport0;
  wire Pre_PE0_Bp0;
  wire Pre_PE0_Bp1;
  wire Pre_PE0_Bp2;
//end pe0 端口定义

//pe1输出端口定义
  reg  [32:0]    PE1_Configure_Inport;
  wire [35:0]    PE1_Outport0;
  wire Pre_PE1_Bp0;
  wire Pre_PE1_Bp1;
  wire Pre_PE1_Bp2;
//end pe1 端口定义

//pe2输出端口定义
  reg  [32:0]    PE2_Configure_Inport;
  wire [35:0]    PE2_Outport0;
  wire Pre_PE2_Bp0;
  wire Pre_PE2_Bp1;
  wire Pre_PE2_Bp2;
//end pe2 端口定义

//pe30输出端口定义
  reg  [32:0]    PE30_Configure_Inport;
  wire [35:0]    PE30_Outport0;
  wire Pre_PE30_Bp0;
  wire Pre_PE30_Bp1;
  wire Pre_PE30_Bp2;
//end pe30 端口定义

//pe3输出端口定义
  reg  [32:0]    PE3_Configure_Inport;
  wire [35:0]    PE3_Outport0;
  wire Pre_PE3_Bp0;
  wire Pre_PE3_Bp1;
  wire Pre_PE3_Bp2;
//end pe3 端口定义

//pe36输出端口定义
  reg  [32:0]    PE36_Configure_Inport;
  wire [35:0]    PE36_Outport0;
  wire Pre_PE36_Bp0;
  wire Pre_PE36_Bp1;
  wire Pre_PE36_Bp2;
//end pe36 端口定义

//pe32输出端口定义
  reg  [32:0]    PE32_Configure_Inport;
  wire [35:0]    PE32_Outport0;
  wire Pre_PE32_Bp0;
  wire Pre_PE32_Bp1;
  wire Pre_PE32_Bp2;
//end pe32 端口定义

//pe5输出端口定义
  reg  [32:0]    PE5_Configure_Inport;
  wire [35:0]    PE5_Outport0;
  wire Pre_PE5_Bp0;
  wire Pre_PE5_Bp1;
  wire Pre_PE5_Bp2;
//end pe5 端口定义

//pe28输出端口定义
  reg  [32:0]    PE28_Configure_Inport;
  wire [35:0]    PE28_Outport0;
  wire Pre_PE28_Bp0;
  wire Pre_PE28_Bp1;
  wire Pre_PE28_Bp2;
//end pe28 端口定义

//pe110输出端口定义
  reg  [32:0]    PE110_Configure_Inport;
  wire [35:0]    PE110_Outport0;
  wire Pre_PE110_Bp0;
  wire Pre_PE110_Bp1;
  wire Pre_PE110_Bp2;
//end pe110 端口定义

//pe6输出端口定义
  reg  [32:0]    PE6_Configure_Inport;
  wire [35:0]    PE6_Outport0;
  wire Pre_PE6_Bp0;
  wire Pre_PE6_Bp1;
  wire Pre_PE6_Bp2;
//end pe6 端口定义

//pe7输出端口定义
  reg  [32:0]    PE7_Configure_Inport;
  wire [35:0]    PE7_Outport0;
  wire Pre_PE7_Bp0;
  wire Pre_PE7_Bp1;
  wire Pre_PE7_Bp2;
//end pe7 端口定义

//pe8输出端口定义
  reg  [32:0]    PE8_Configure_Inport;
  wire [35:0]    PE8_Outport0;
  wire Pre_PE8_Bp0;
  wire Pre_PE8_Bp1;
  wire Pre_PE8_Bp2;
//end pe8 端口定义

//pe9输出端口定义
  reg  [32:0]    PE9_Configure_Inport;
  wire [35:0]    PE9_Outport0;
  wire Pre_PE9_Bp0;
  wire Pre_PE9_Bp1;
  wire Pre_PE9_Bp2;
//end pe9 端口定义

//pe29输出端口定义
  reg  [32:0]    PE29_Configure_Inport;
  wire [35:0]    PE29_Outport0;
  wire Pre_PE29_Bp0;
  wire Pre_PE29_Bp1;
  wire Pre_PE29_Bp2;
//end pe29 端口定义

//pe31输出端口定义
  reg  [32:0]    PE31_Configure_Inport;
  wire [35:0]    PE31_Outport0;
  wire Pre_PE31_Bp0;
  wire Pre_PE31_Bp1;
  wire Pre_PE31_Bp2;
//end pe31 端口定义

//pe10输出端口定义
  reg  [32:0]    PE10_Configure_Inport;
  wire [35:0]    PE10_Outport0;
  wire Pre_PE10_Bp0;
  wire Pre_PE10_Bp1;
  wire Pre_PE10_Bp2;
//end pe10 端口定义

//pe37输出端口定义
  reg  [32:0]    PE37_Configure_Inport;
  wire [35:0]    PE37_Outport0;
  wire Pre_PE37_Bp0;
  wire Pre_PE37_Bp1;
  wire Pre_PE37_Bp2;
//end pe37 端口定义

//pe11输出端口定义
  reg  [32:0]    PE11_Configure_Inport;
  wire [35:0]    PE11_Outport0;
  wire Pre_PE11_Bp0;
  wire Pre_PE11_Bp1;
  wire Pre_PE11_Bp2;
//end pe11 端口定义

//pe12输出端口定义
  reg  [32:0]    PE12_Configure_Inport;
  wire [35:0]    PE12_Outport0;
  wire Pre_PE12_Bp0;
  wire Pre_PE12_Bp1;
  wire Pre_PE12_Bp2;
//end pe12 端口定义

//pe13输出端口定义
  reg  [32:0]    PE13_Configure_Inport;
  wire [35:0]    PE13_Outport0;
  wire Pre_PE13_Bp0;
  wire Pre_PE13_Bp1;
  wire Pre_PE13_Bp2;
//end pe13 端口定义

//pe109输出端口定义
  reg  [32:0]    PE109_Configure_Inport;
  wire [35:0]    PE109_Outport0;
  wire Pre_PE109_Bp0;
  wire Pre_PE109_Bp1;
  wire Pre_PE109_Bp2;
//end pe109 端口定义

//pe100输出端口定义
  reg  [32:0]    PE100_Configure_Inport;
  wire [35:0]    PE100_Outport0;
  wire Pre_PE100_Bp0;
  wire Pre_PE100_Bp1;
  wire Pre_PE100_Bp2;
//end pe100 端口定义

//pe102输出端口定义
  reg  [32:0]    PE102_Configure_Inport;
  wire [35:0]    PE102_Outport0;
  wire Pre_PE102_Bp0;
  wire Pre_PE102_Bp1;
  wire Pre_PE102_Bp2;
//end pe102 端口定义

//pe103输出端口定义
  reg  [32:0]    PE103_Configure_Inport;
  wire [35:0]    PE103_Outport0;
  wire Pre_PE103_Bp0;
  wire Pre_PE103_Bp1;
  wire Pre_PE103_Bp2;
//end pe103 端口定义

//pe104输出端口定义
  reg  [32:0]    PE104_Configure_Inport;
  wire [35:0]    PE104_Outport0;
  wire Pre_PE104_Bp0;
  wire Pre_PE104_Bp1;
  wire Pre_PE104_Bp2;
//end pe104 端口定义

//pe14输出端口定义
  reg  [32:0]    PE14_Configure_Inport;
  wire [35:0]    PE14_Outport0;
  wire Pre_PE14_Bp0;
  wire Pre_PE14_Bp1;
  wire Pre_PE14_Bp2;
//end pe14 端口定义

//pe21输出端口定义
  reg  [32:0]    PE21_Configure_Inport;
  wire [35:0]    PE21_Outport0;
  wire Pre_PE21_Bp0;
  wire Pre_PE21_Bp1;
  wire Pre_PE21_Bp2;
//end pe21 端口定义

//pe15输出端口定义
  reg  [32:0]    PE15_Configure_Inport;
  wire [35:0]    PE15_Outport0;
  wire Pre_PE15_Bp0;
  wire Pre_PE15_Bp1;
  wire Pre_PE15_Bp2;
//end pe15 端口定义

//pe16输出端口定义
  reg  [32:0]    PE16_Configure_Inport;
  wire [35:0]    PE16_Outport0;
  wire Pre_PE16_Bp0;
  wire Pre_PE16_Bp1;
  wire Pre_PE16_Bp2;
//end pe16 端口定义

//pe17输出端口定义
  reg  [32:0]    PE17_Configure_Inport;
  wire [35:0]    PE17_Outport0;
  wire Pre_PE17_Bp0;
  wire Pre_PE17_Bp1;
  wire Pre_PE17_Bp2;
//end pe17 端口定义

//pe101输出端口定义
  reg  [32:0]    PE101_Configure_Inport;
  wire [35:0]    PE101_Outport0;
  wire Pre_PE101_Bp0;
  wire Pre_PE101_Bp1;
  wire Pre_PE101_Bp2;
//end pe101 端口定义

//pe19输出端口定义
  reg  [32:0]    PE19_Configure_Inport;
  wire [35:0]    PE19_Outport0;
  wire Pre_PE19_Bp0;
  wire Pre_PE19_Bp1;
  wire Pre_PE19_Bp2;
//end pe19 端口定义

//pe22输出端口定义
  reg  [32:0]    PE22_Configure_Inport;
  wire [35:0]    PE22_Outport0;
  wire Pre_PE22_Bp0;
  wire Pre_PE22_Bp1;
  wire Pre_PE22_Bp2;
//end pe22 端口定义

//pe23输出端口定义
  reg  [32:0]    PE23_Configure_Inport;
  wire [35:0]    PE23_Outport0;
  wire Pre_PE23_Bp0;
  wire Pre_PE23_Bp1;
  wire Pre_PE23_Bp2;
//end pe23 端口定义

//pe24输出端口定义
  reg  [32:0]    PE24_Configure_Inport;
  wire [35:0]    PE24_Outport0;
  wire Pre_PE24_Bp0;
  wire Pre_PE24_Bp1;
  wire Pre_PE24_Bp2;
//end pe24 端口定义

//pe111输出端口定义
  reg  [32:0]    PE111_Configure_Inport;
  wire [35:0]    PE111_Outport0;
  wire Pre_PE111_Bp0;
  wire Pre_PE111_Bp1;
  wire Pre_PE111_Bp2;
//end pe111 端口定义

//pe26输出端口定义
  reg  [32:0]    PE26_Configure_Inport;
  wire [35:0]    PE26_Outport0;
  wire Pre_PE26_Bp0;
  wire Pre_PE26_Bp1;
  wire Pre_PE26_Bp2;
//end pe26 端口定义

//pe27输出端口定义
  reg  [32:0]    PE27_Configure_Inport;
  wire [35:0]    PE27_Outport0;
  wire Pre_PE27_Bp0;
  wire Pre_PE27_Bp1;
  wire Pre_PE27_Bp2;
//end pe27 端口定义

//pe25输出端口定义
  reg  [32:0]    PE25_Configure_Inport;
  wire [35:0]    PE25_Outport0;
  wire Pre_PE25_Bp0;
  wire Pre_PE25_Bp1;
  wire Pre_PE25_Bp2;
//end pe25 端口定义

//pe38例化
PE_top  pe38_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(36'b0),
    .PE_Inport1(PE38_Inport1),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE0_Bp0),
    .Post_PE_Bp1(Pre_PE1_Bp0),
    .Post_PE_Bp2(Pre_PE2_Bp0),
    .Post_PE_Bp3(Pre_PE5_Bp1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE38_Configure_Inport),
    .PE_Outport0(PE38_Outport0),
    .Pre_PE_Bp0(Pre_PE38_Bp0),
    .Pre_PE_Bp1(Pre_PE38_Bp1),
    .Pre_PE_Bp2(Pre_PE38_Bp2)
);
//end pe38 例化
    
//pe0例化
PE_top  pe0_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE38_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE2_Bp2),
    .Post_PE_Bp1(Pre_PE30_Bp1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE0_Configure_Inport),
    .PE_Outport0(PE0_Outport0),
    .Pre_PE_Bp0(Pre_PE0_Bp0),
    .Pre_PE_Bp1(Pre_PE0_Bp1),
    .Pre_PE_Bp2(Pre_PE0_Bp2)
);
//end pe0 例化
    
//pe1例化
PE_top  pe1_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE38_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE3_Bp0),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE1_Configure_Inport),
    .PE_Outport0(PE1_Outport0),
    .Pre_PE_Bp0(Pre_PE1_Bp0),
    .Pre_PE_Bp1(Pre_PE1_Bp1),
    .Pre_PE_Bp2(Pre_PE1_Bp2)
);
//end pe1 例化
    
//pe2例化
PE_top  pe2_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE38_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(PE0_Outport0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE36_Bp2),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE2_Configure_Inport),
    .PE_Outport0(PE2_Outport0),
    .Pre_PE_Bp0(Pre_PE2_Bp0),
    .Pre_PE_Bp1(Pre_PE2_Bp1),
    .Pre_PE_Bp2(Pre_PE2_Bp2)
);
//end pe2 例化
    
//pe30例化
PE_top  pe30_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(36'b0),
    .PE_Inport1(PE0_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE3_Bp2),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE30_Configure_Inport),
    .PE_Outport0(PE30_Outport0),
    .Pre_PE_Bp0(Pre_PE30_Bp0),
    .Pre_PE_Bp1(Pre_PE30_Bp1),
    .Pre_PE_Bp2(Pre_PE30_Bp2)
);
//end pe30 例化
    
//pe3例化
PE_top  pe3_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE1_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(PE30_Outport0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE36_Bp1),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE3_Configure_Inport),
    .PE_Outport0(PE3_Outport0),
    .Pre_PE_Bp0(Pre_PE3_Bp0),
    .Pre_PE_Bp1(Pre_PE3_Bp1),
    .Pre_PE_Bp2(Pre_PE3_Bp2)
);
//end pe3 例化
    
//pe36例化
PE_top  pe36_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(36'b0),
    .PE_Inport1(PE3_Outport0),
    .PE_Inport2(PE2_Outport0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE32_Bp1),
    .Post_PE_Bp1(Pre_PE110_Bp1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE36_Configure_Inport),
    .PE_Outport0(PE36_Outport0),
    .Pre_PE_Bp0(Pre_PE36_Bp0),
    .Pre_PE_Bp1(Pre_PE36_Bp1),
    .Pre_PE_Bp2(Pre_PE36_Bp2)
);
//end pe36 例化
    
//pe32例化
PE_top  pe32_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(36'b0),
    .PE_Inport1(PE36_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE5_Bp0),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE32_Configure_Inport),
    .PE_Outport0(PE32_Outport0),
    .Pre_PE_Bp0(Pre_PE32_Bp0),
    .Pre_PE_Bp1(Pre_PE32_Bp1),
    .Pre_PE_Bp2(Pre_PE32_Bp2)
);
//end pe32 例化
    
//pe5例化
PE_top  pe5_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE32_Outport0),
    .PE_Inport1(PE38_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE28_Bp0),
    .Post_PE_Bp1(Pre_PE9_Bp0),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE5_Configure_Inport),
    .PE_Outport0(PE5_Outport0),
    .Pre_PE_Bp0(Pre_PE5_Bp0),
    .Pre_PE_Bp1(Pre_PE5_Bp1),
    .Pre_PE_Bp2(Pre_PE5_Bp2)
);
//end pe5 例化
    
//pe28例化
PE_top  pe28_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE5_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE13_Bp0),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE28_Configure_Inport),
    .PE_Outport0(PE28_Outport0),
    .Pre_PE_Bp0(Pre_PE28_Bp0),
    .Pre_PE_Bp1(Pre_PE28_Bp1),
    .Pre_PE_Bp2(Pre_PE28_Bp2)
);
//end pe28 例化
    
//pe110例化
PE_top  pe110_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(36'b0),
    .PE_Inport1(PE36_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE6_Bp0),
    .Post_PE_Bp1(Pre_PE8_Bp0),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE110_Configure_Inport),
    .PE_Outport0(PE110_Outport0),
    .Pre_PE_Bp0(Pre_PE110_Bp0),
    .Pre_PE_Bp1(Pre_PE110_Bp1),
    .Pre_PE_Bp2(Pre_PE110_Bp2)
);
//end pe110 例化
    
//pe6例化
PE_top  pe6_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE110_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE7_Bp0),
    .Post_PE_Bp1(Pre_PE31_Bp0),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE6_Configure_Inport),
    .PE_Outport0(PE6_Outport0),
    .Pre_PE_Bp0(Pre_PE6_Bp0),
    .Pre_PE_Bp1(Pre_PE6_Bp1),
    .Pre_PE_Bp2(Pre_PE6_Bp2)
);
//end pe6 例化
    
//pe7例化
PE_top  pe7_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE6_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE10_Bp1),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE7_Configure_Inport),
    .PE_Outport0(PE7_Outport0),
    .Pre_PE_Bp0(Pre_PE7_Bp0),
    .Pre_PE_Bp1(Pre_PE7_Bp1),
    .Pre_PE_Bp2(Pre_PE7_Bp2)
);
//end pe7 例化
    
//pe8例化
PE_top  pe8_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE110_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE12_Bp1),
    .Post_PE_Bp1(Pre_PE13_Bp1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE8_Configure_Inport),
    .PE_Outport0(PE8_Outport0),
    .Pre_PE_Bp0(Pre_PE8_Bp0),
    .Pre_PE_Bp1(Pre_PE8_Bp1),
    .Pre_PE_Bp2(Pre_PE8_Bp2)
);
//end pe8 例化
    
//pe9例化
PE_top  pe9_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE5_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE29_Bp0),
    .Post_PE_Bp1(Pre_PE109_Bp1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE9_Configure_Inport),
    .PE_Outport0(PE9_Outport0),
    .Pre_PE_Bp0(Pre_PE9_Bp0),
    .Pre_PE_Bp1(Pre_PE9_Bp1),
    .Pre_PE_Bp2(Pre_PE9_Bp2)
);
//end pe9 例化
    
//pe29例化
PE_top  pe29_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE9_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE10_Bp0),
    .Post_PE_Bp1(Pre_PE12_Bp0),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE29_Configure_Inport),
    .PE_Outport0(PE29_Outport0),
    .Pre_PE_Bp0(Pre_PE29_Bp0),
    .Pre_PE_Bp1(Pre_PE29_Bp1),
    .Pre_PE_Bp2(Pre_PE29_Bp2)
);
//end pe29 例化
    
//pe31例化
PE_top  pe31_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE6_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE100_Bp1),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE31_Configure_Inport),
    .PE_Outport0(PE31_Outport0),
    .Pre_PE_Bp0(Pre_PE31_Bp0),
    .Pre_PE_Bp1(Pre_PE31_Bp1),
    .Pre_PE_Bp2(Pre_PE31_Bp2)
);
//end pe31 例化
    
//pe10例化
PE_top  pe10_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE29_Outport0),
    .PE_Inport1(PE7_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE37_Bp0),
    .Post_PE_Bp1(Pre_PE11_Bp0),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE10_Configure_Inport),
    .PE_Outport0(PE10_Outport0),
    .Pre_PE_Bp0(Pre_PE10_Bp0),
    .Pre_PE_Bp1(Pre_PE10_Bp1),
    .Pre_PE_Bp2(Pre_PE10_Bp2)
);
//end pe10 例化
    
//pe37例化
PE_top  pe37_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE10_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE102_Bp1),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE37_Configure_Inport),
    .PE_Outport0(PE37_Outport0),
    .Pre_PE_Bp0(Pre_PE37_Bp0),
    .Pre_PE_Bp1(Pre_PE37_Bp1),
    .Pre_PE_Bp2(Pre_PE37_Bp2)
);
//end pe37 例化
    
//pe11例化
PE_top  pe11_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE10_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE103_Bp1),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE11_Configure_Inport),
    .PE_Outport0(PE11_Outport0),
    .Pre_PE_Bp0(Pre_PE11_Bp0),
    .Pre_PE_Bp1(Pre_PE11_Bp1),
    .Pre_PE_Bp2(Pre_PE11_Bp2)
);
//end pe11 例化
    
//pe12例化
PE_top  pe12_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE29_Outport0),
    .PE_Inport1(PE8_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE104_Bp1),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE12_Configure_Inport),
    .PE_Outport0(PE12_Outport0),
    .Pre_PE_Bp0(Pre_PE12_Bp0),
    .Pre_PE_Bp1(Pre_PE12_Bp1),
    .Pre_PE_Bp2(Pre_PE12_Bp2)
);
//end pe12 例化
    
//pe13例化
PE_top  pe13_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE28_Outport0),
    .PE_Inport1(PE8_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE101_Bp1),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE13_Configure_Inport),
    .PE_Outport0(PE13_Outport0),
    .Pre_PE_Bp0(Pre_PE13_Bp0),
    .Pre_PE_Bp1(Pre_PE13_Bp1),
    .Pre_PE_Bp2(Pre_PE13_Bp2)
);
//end pe13 例化
    
//pe109例化
PE_top  pe109_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(36'b0),
    .PE_Inport1(PE9_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE14_Bp1),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE109_Configure_Inport),
    .PE_Outport0(PE109_Outport0),
    .Pre_PE_Bp0(Pre_PE109_Bp0),
    .Pre_PE_Bp1(Pre_PE109_Bp1),
    .Pre_PE_Bp2(Pre_PE109_Bp2)
);
//end pe109 例化
    
//pe100例化
PE_top  pe100_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(36'b0),
    .PE_Inport1(PE31_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE14_Bp0),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE100_Configure_Inport),
    .PE_Outport0(PE100_Outport0),
    .Pre_PE_Bp0(Pre_PE100_Bp0),
    .Pre_PE_Bp1(Pre_PE100_Bp1),
    .Pre_PE_Bp2(Pre_PE100_Bp2)
);
//end pe100 例化
    
//pe102例化
PE_top  pe102_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(36'b0),
    .PE_Inport1(PE37_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE15_Bp0),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE102_Configure_Inport),
    .PE_Outport0(PE102_Outport0),
    .Pre_PE_Bp0(Pre_PE102_Bp0),
    .Pre_PE_Bp1(Pre_PE102_Bp1),
    .Pre_PE_Bp2(Pre_PE102_Bp2)
);
//end pe102 例化
    
//pe103例化
PE_top  pe103_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(36'b0),
    .PE_Inport1(PE11_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE16_Bp0),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE103_Configure_Inport),
    .PE_Outport0(PE103_Outport0),
    .Pre_PE_Bp0(Pre_PE103_Bp0),
    .Pre_PE_Bp1(Pre_PE103_Bp1),
    .Pre_PE_Bp2(Pre_PE103_Bp2)
);
//end pe103 例化
    
//pe104例化
PE_top  pe104_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(36'b0),
    .PE_Inport1(PE12_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE17_Bp0),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE104_Configure_Inport),
    .PE_Outport0(PE104_Outport0),
    .Pre_PE_Bp0(Pre_PE104_Bp0),
    .Pre_PE_Bp1(Pre_PE104_Bp1),
    .Pre_PE_Bp2(Pre_PE104_Bp2)
);
//end pe104 例化
    
//pe14例化
PE_top  pe14_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE100_Outport0),
    .PE_Inport1(PE109_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE21_Bp2),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE14_Configure_Inport),
    .PE_Outport0(PE14_Outport0),
    .Pre_PE_Bp0(Pre_PE14_Bp0),
    .Pre_PE_Bp1(Pre_PE14_Bp1),
    .Pre_PE_Bp2(Pre_PE14_Bp2)
);
//end pe14 例化
    
//pe21例化
PE_top  pe21_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(36'b0),
    .PE_Inport1(36'b0),
    .PE_Inport2(PE14_Outport0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE15_Bp1),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE21_Configure_Inport),
    .PE_Outport0(PE21_Outport0),
    .Pre_PE_Bp0(Pre_PE21_Bp0),
    .Pre_PE_Bp1(Pre_PE21_Bp1),
    .Pre_PE_Bp2(Pre_PE21_Bp2)
);
//end pe21 例化
    
//pe15例化
PE_top  pe15_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE102_Outport0),
    .PE_Inport1(PE21_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE111_Bp1),
    .Post_PE_Bp1(Pre_PE27_Bp1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE15_Configure_Inport),
    .PE_Outport0(PE15_Outport0),
    .Pre_PE_Bp0(Pre_PE15_Bp0),
    .Pre_PE_Bp1(Pre_PE15_Bp1),
    .Pre_PE_Bp2(Pre_PE15_Bp2)
);
//end pe15 例化
    
//pe16例化
PE_top  pe16_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE103_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE22_Bp1),
    .Post_PE_Bp1(Pre_PE24_Bp0),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE16_Configure_Inport),
    .PE_Outport0(PE16_Outport0),
    .Pre_PE_Bp0(Pre_PE16_Bp0),
    .Pre_PE_Bp1(Pre_PE16_Bp1),
    .Pre_PE_Bp2(Pre_PE16_Bp2)
);
//end pe16 例化
    
//pe17例化
PE_top  pe17_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE104_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE22_Bp0),
    .Post_PE_Bp1(Pre_PE24_Bp1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE17_Configure_Inport),
    .PE_Outport0(PE17_Outport0),
    .Pre_PE_Bp0(Pre_PE17_Bp0),
    .Pre_PE_Bp1(Pre_PE17_Bp1),
    .Pre_PE_Bp2(Pre_PE17_Bp2)
);
//end pe17 例化
    
//pe101例化
PE_top  pe101_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(36'b0),
    .PE_Inport1(PE13_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE19_Bp0),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE101_Configure_Inport),
    .PE_Outport0(PE101_Outport0),
    .Pre_PE_Bp0(Pre_PE101_Bp0),
    .Pre_PE_Bp1(Pre_PE101_Bp1),
    .Pre_PE_Bp2(Pre_PE101_Bp2)
);
//end pe101 例化
    
//pe19例化
PE_top  pe19_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE101_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(1'b1),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE19_Configure_Inport),
    .PE_Outport0(PE19_Outport0),
    .Pre_PE_Bp0(Pre_PE19_Bp0),
    .Pre_PE_Bp1(Pre_PE19_Bp1),
    .Pre_PE_Bp2(Pre_PE19_Bp2)
);
//end pe19 例化
    
//pe22例化
PE_top  pe22_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE17_Outport0),
    .PE_Inport1(PE16_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE23_Bp2),
    .Post_PE_Bp1(Pre_PE24_Bp2),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE22_Configure_Inport),
    .PE_Outport0(PE22_Outport0),
    .Pre_PE_Bp0(Pre_PE22_Bp0),
    .Pre_PE_Bp1(Pre_PE22_Bp1),
    .Pre_PE_Bp2(Pre_PE22_Bp2)
);
//end pe22 例化
    
//pe23例化
PE_top  pe23_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(36'b0),
    .PE_Inport1(36'b0),
    .PE_Inport2(PE22_Outport0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE25_Bp0),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE23_Configure_Inport),
    .PE_Outport0(PE23_Outport0),
    .Pre_PE_Bp0(Pre_PE23_Bp0),
    .Pre_PE_Bp1(Pre_PE23_Bp1),
    .Pre_PE_Bp2(Pre_PE23_Bp2)
);
//end pe23 例化
    
//pe24例化
PE_top  pe24_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE16_Outport0),
    .PE_Inport1(PE17_Outport0),
    .PE_Inport2(PE22_Outport0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE26_Bp1),
    .Post_PE_Bp1(Pre_PE27_Bp0),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE24_Configure_Inport),
    .PE_Outport0(PE24_Outport0),
    .Pre_PE_Bp0(Pre_PE24_Bp0),
    .Pre_PE_Bp1(Pre_PE24_Bp1),
    .Pre_PE_Bp2(Pre_PE24_Bp2)
);
//end pe24 例化
    
//pe111例化
PE_top  pe111_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(36'b0),
    .PE_Inport1(PE15_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE26_Bp0),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE111_Configure_Inport),
    .PE_Outport0(PE111_Outport0),
    .Pre_PE_Bp0(Pre_PE111_Bp0),
    .Pre_PE_Bp1(Pre_PE111_Bp1),
    .Pre_PE_Bp2(Pre_PE111_Bp2)
);
//end pe111 例化
    
//pe26例化
PE_top  pe26_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE111_Outport0),
    .PE_Inport1(PE24_Outport0),
    .PE_Inport2(36'b0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(Pre_PE27_Bp2),
    .Post_PE_Bp1(Pre_PE25_Bp2),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE26_Configure_Inport),
    .PE_Outport0(PE26_Outport0),
    .Pre_PE_Bp0(Pre_PE26_Bp0),
    .Pre_PE_Bp1(Pre_PE26_Bp1),
    .Pre_PE_Bp2(Pre_PE26_Bp2)
);
//end pe26 例化
    
//pe27例化
PE_top  pe27_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE24_Outport0),
    .PE_Inport1(PE15_Outport0),
    .PE_Inport2(PE26_Outport0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(1'b1),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE27_Configure_Inport),
    .PE_Outport0(PE27_Outport0),
    .Pre_PE_Bp0(Pre_PE27_Bp0),
    .Pre_PE_Bp1(Pre_PE27_Bp1),
    .Pre_PE_Bp2(Pre_PE27_Bp2)
);
//end pe27 例化
    
//pe25例化
PE_top  pe25_top(
    .clk(clk),
    .reset(rst),
    .PE_Inport0(PE23_Outport0),
    .PE_Inport1(36'b0),
    .PE_Inport2(PE26_Outport0),
    .PE_Bus_Port0(4'b0),
    .Post_PE_Bp0(1'b1),
    .Post_PE_Bp1(1'b1),
    .Post_PE_Bp2(1'b1),
    .Post_PE_Bp3(1'b1),
    .Post_PE_Bp4(1'b1),
    .Post_PE_Bp5(1'b1),
    .Post_PE_Bp6(1'b1),
    .Post_PE_Bp7(1'b1),
    .PE_Configure_Inport(PE25_Configure_Inport),
    .PE_Outport0(PE25_Outport0),
    .Pre_PE_Bp0(Pre_PE25_Bp0),
    .Pre_PE_Bp1(Pre_PE25_Bp1),
    .Pre_PE_Bp2(Pre_PE25_Bp2)
);
//end pe25 例化
    
  initial begin
    rst <=1'b1;
    clk <=1'b0;
    PE38_Configure_Inport <={1'b1,7'b000_0000,3'b101,1'b1,5'd5,3'b101,4'b0100,2'b01,1'd0,4'd2,2'd0};
    PE0_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd5,3'b010,4'b1000,2'b00,1'd0,4'd0,2'd0};
    PE1_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd4,3'b010,4'b1000,2'b00,1'd0,4'd0,2'd0};
    PE2_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd13,3'b010,4'b1001,2'b00,1'd0,4'd0,2'd0};
    PE30_Configure_Inport <={1'b1,7'b000_0000,3'b000,1'b1,5'd18,3'b000,4'b0010,2'b00,1'd0,4'd0,2'd0};
    PE3_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd13,3'b010,4'b1001,2'b00,1'd0,4'd0,2'd0};
    PE36_Configure_Inport <={1'b1,7'b000_0000,3'b100,1'b1,5'd5,3'b101,4'b0101,2'b01,1'd0,4'd10,2'd0};
    PE32_Configure_Inport <={1'b1,7'b000_0000,3'b100,1'b1,5'd4,3'b100,4'b0010,2'b00,1'd0,4'd0,2'd0};
    PE5_Configure_Inport <={1'b1,7'b000_0000,3'b000,1'b1,5'd3,3'b010,4'b1010,2'b00,1'd0,4'd0,2'd0};
    PE28_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd3,3'b010,4'b1000,2'b00,1'd0,4'd0,2'd0};
    PE110_Configure_Inport <={1'b1,7'b000_0000,3'b100,1'b1,5'd3,3'b100,4'b0010,2'b00,1'd0,4'd0,2'd0};
    PE6_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd4,3'b010,4'b1000,2'b00,1'd0,4'd0,2'd0};
    PE7_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd2,3'b010,4'b1000,2'b00,1'd0,4'd0,2'd0};
    PE8_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd2,3'b010,4'b1000,2'b00,1'd0,4'd0,2'd0};
    PE9_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd4,3'b010,4'b1000,2'b00,1'd0,4'd0,2'd0};
    PE29_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd3,3'b010,4'b1000,2'b00,1'd0,4'd0,2'd0};
    PE31_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd3,3'b010,4'b1000,2'b00,1'd0,4'd0,2'd0};
    PE10_Configure_Inport <={1'b1,7'b000_0000,3'b000,1'b1,5'd3,3'b000,4'b1010,2'b00,1'd0,4'd0,2'd0};
    PE37_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd3,3'b010,4'b1000,2'b00,1'd0,4'd0,2'd0};
    PE11_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd3,3'b010,4'b1000,2'b00,1'd0,4'd0,2'd0};
    PE12_Configure_Inport <={1'b1,7'b000_0000,3'b000,1'b1,5'd3,3'b000,4'b1010,2'b00,1'd0,4'd0,2'd0};
    PE13_Configure_Inport <={1'b1,7'b000_0000,3'b000,1'b1,5'd3,3'b000,4'b1010,2'b00,1'd0,4'd0,2'd0};
    PE109_Configure_Inport <={1'b1,7'b000_0000,3'b100,1'b1,5'd3,3'b100,4'b0010,2'b00,1'd0,4'd0,2'd0};
    PE100_Configure_Inport <={1'b1,7'b000_0000,3'b100,1'b1,5'd3,3'b100,4'b0010,2'b00,1'd0,4'd0,2'd0};
    PE102_Configure_Inport <={1'b1,7'b000_0000,3'b100,1'b1,5'd3,3'b100,4'b0010,2'b00,1'd0,4'd0,2'd0};
    PE103_Configure_Inport <={1'b1,7'b000_0000,3'b100,1'b1,5'd3,3'b100,4'b0010,2'b00,1'd0,4'd0,2'd0};
    PE104_Configure_Inport <={1'b1,7'b000_0000,3'b100,1'b1,5'd3,3'b100,4'b0010,2'b00,1'd0,4'd0,2'd0};
    PE14_Configure_Inport <={1'b1,7'b000_0000,3'b000,1'b1,5'd7,3'b000,4'b1010,2'b00,1'd0,4'd0,2'd0};
    PE21_Configure_Inport <={1'b1,7'b000_0000,3'b110,1'b1,5'd13,3'b110,4'b0001,2'b00,1'd0,4'd0,2'd0};
    PE15_Configure_Inport <={1'b1,7'b000_0000,3'b000,1'b1,5'd3,3'b000,4'b1010,2'b00,1'd0,4'd0,2'd0};
    PE16_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd4,3'b010,4'b1000,2'b00,1'd0,4'd0,2'd0};
    PE17_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd4,3'b010,4'b1000,2'b00,1'd0,4'd0,2'd0};
    PE101_Configure_Inport <={1'b1,7'b000_0000,3'b100,1'b1,5'd3,3'b100,4'b0010,2'b00,1'd0,4'd0,2'd0};
    PE19_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd3,3'b010,4'b1000,2'b00,1'd0,4'd0,2'd0};
    PE22_Configure_Inport <={1'b1,7'b000_0000,3'b000,1'b1,5'd5,3'b000,4'b1010,2'b00,1'd0,4'd0,2'd0};
    PE23_Configure_Inport <={1'b1,7'b000_0000,3'b110,1'b1,5'd13,3'b110,4'b0001,2'b00,1'd0,4'd0,2'd0};
    PE24_Configure_Inport <={1'b1,7'b000_0000,3'b000,1'b1,5'd13,3'b000,4'b1011,2'b00,1'd0,4'd0,2'd0};
    PE111_Configure_Inport <={1'b1,7'b000_0000,3'b100,1'b1,5'd3,3'b100,4'b0010,2'b00,1'd0,4'd0,2'd0};
    PE26_Configure_Inport <={1'b1,7'b000_0000,3'b000,1'b1,5'd5,3'b000,4'b1010,2'b00,1'd0,4'd0,2'd0};
    PE27_Configure_Inport <={1'b1,7'b000_0000,3'b000,1'b1,5'd13,3'b000,4'b1011,2'b00,1'd0,4'd0,2'd0};
    PE25_Configure_Inport <={1'b1,7'b000_0000,3'b010,1'b1,5'd13,3'b010,4'b1001,2'b00,1'd0,4'd0,2'd0};
    #2 rst <= ~rst;
    #1 rst <= ~rst;
    #10 PE30_Configure_Inport <=33'd0;
        PE102_Configure_Inport <={1'b1,32'd0};
        PE38_Configure_Inport <={1'b1,32'd2};
        PE32_Configure_Inport <={1'b1,32'd0};
        PE0_Configure_Inport <={1'b1,32'd65};
        PE1_Configure_Inport <={1'b1,32'd64};
        PE2_Configure_Inport <={1'b1,32'd65};
        PE3_Configure_Inport <={1'b1,32'd1};
        PE100_Configure_Inport <={1'b1,32'd0};
        PE36_Configure_Inport <={1'b1,32'd1};
        PE5_Configure_Inport <=33'd0;
        PE28_Configure_Inport <={1'b1,32'd144};
        PE110_Configure_Inport <={1'b1,32'd0};
        PE6_Configure_Inport <={1'b1,32'd1};
        PE7_Configure_Inport <={1'b1,32'd72};
        PE8_Configure_Inport <={1'b1,32'd72};
        PE9_Configure_Inport <={1'b1,32'd1};
        PE29_Configure_Inport <={1'b1,32'd144};
        PE31_Configure_Inport <={1'b1,32'd72};
        PE10_Configure_Inport <=33'd0;
        PE101_Configure_Inport <={1'b1,32'd0};
        PE37_Configure_Inport <={1'b1,32'd0};
        PE11_Configure_Inport <={1'b1,32'd1};
        PE12_Configure_Inport <=33'd0;
        PE13_Configure_Inport <=33'd0;
        PE109_Configure_Inport <={1'b1,32'd0};
        PE103_Configure_Inport <={1'b1,32'd0};
        PE104_Configure_Inport <={1'b1,32'd0};
        PE14_Configure_Inport <=33'd0;
        PE21_Configure_Inport <={1'b1,32'd1};
        PE15_Configure_Inport <=33'd0;
        PE16_Configure_Inport <={1'b1,32'd1};
        PE17_Configure_Inport <={1'b1,32'd1};
        PE19_Configure_Inport <={1'b1,32'd9288};
        PE22_Configure_Inport <=33'd0;
        PE23_Configure_Inport <={1'b1,32'd94};
        PE24_Configure_Inport <=33'd0;
        PE111_Configure_Inport <={1'b1,32'd0};
        PE26_Configure_Inport <=33'd0;
        PE27_Configure_Inport <=33'd0;
        PE25_Configure_Inport <={1'b1,32'd47};
    #10 PE102_Configure_Inport <=33'd0;
        PE38_Configure_Inport <={1'b1,32'd129};
        PE32_Configure_Inport <=33'd0;
        PE0_Configure_Inport <=33'd0;
        PE1_Configure_Inport <=33'd0;
        PE2_Configure_Inport <=33'd0;
        PE3_Configure_Inport <=33'd0;
        PE100_Configure_Inport <=33'd0;
        PE36_Configure_Inport <=33'd0;
        PE28_Configure_Inport <=33'd0;
        PE110_Configure_Inport <=33'd0;
        PE6_Configure_Inport <=33'd0;
        PE7_Configure_Inport <=33'd0;
        PE8_Configure_Inport <=33'd0;
        PE9_Configure_Inport <=33'd0;
        PE29_Configure_Inport <=33'd0;
        PE31_Configure_Inport <=33'd0;
        PE101_Configure_Inport <=33'd0;
        PE37_Configure_Inport <=33'd0;
        PE11_Configure_Inport <=33'd0;
        PE109_Configure_Inport <=33'd0;
        PE103_Configure_Inport <=33'd0;
        PE104_Configure_Inport <=33'd0;
        PE21_Configure_Inport <={1'b1,32'd-1};
        PE16_Configure_Inport <=33'd0;
        PE17_Configure_Inport <=33'd0;
        PE19_Configure_Inport <=33'd0;
        PE23_Configure_Inport <={1'b1,32'd60};
        PE111_Configure_Inport <=33'd0;
        PE25_Configure_Inport <=33'd0;
    #10 PE38_Configure_Inport <=33'd0;
        PE21_Configure_Inport <=33'd0;
        PE23_Configure_Inport <=33'd0;
    #10 PE38_Inport1 <= {4'b1100,32'd0};
    #10 PE38_Inport1 <= {4'b0000,32'd0};
  end
  initial begin
      filez=$fopen("./data_flow_rtl","w");
        for(i=0;i<100;i=i+1) begin
            @(posedge clk);
            #1
            if(PE38_Outport0[35:33]!=3'b000&&PE38_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE38.vbl=%b,value=%d@clk %d\n",PE38_Outport0[35:33],PE38_Outport0[31:0],i);
            end
            if(PE0_Outport0[35:33]!=3'b000&&PE0_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE0.vbl=%b,value=%d@clk %d\n",PE0_Outport0[35:33],PE0_Outport0[31:0],i);
            end
            if(PE1_Outport0[35:33]!=3'b000&&PE1_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE1.vbl=%b,value=%d@clk %d\n",PE1_Outport0[35:33],PE1_Outport0[31:0],i);
            end
            if(PE2_Outport0[35:33]!=3'b000&&PE2_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE2.vbl=%b,value=%d@clk %d\n",PE2_Outport0[35:33],PE2_Outport0[31:0],i);
            end
            if(PE30_Outport0[35:33]!=3'b000&&PE30_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE30.vbl=%b,value=%d@clk %d\n",PE30_Outport0[35:33],PE30_Outport0[31:0],i);
            end
            if(PE3_Outport0[35:33]!=3'b000&&PE3_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE3.vbl=%b,value=%d@clk %d\n",PE3_Outport0[35:33],PE3_Outport0[31:0],i);
            end
            if(PE36_Outport0[35:33]!=3'b000&&PE36_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE36.vbl=%b,value=%d@clk %d\n",PE36_Outport0[35:33],PE36_Outport0[31:0],i);
            end
            if(PE32_Outport0[35:33]!=3'b000&&PE32_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE32.vbl=%b,value=%d@clk %d\n",PE32_Outport0[35:33],PE32_Outport0[31:0],i);
            end
            if(PE5_Outport0[35:33]!=3'b000&&PE5_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE5.vbl=%b,value=%d@clk %d\n",PE5_Outport0[35:33],PE5_Outport0[31:0],i);
            end
            if(PE28_Outport0[35:33]!=3'b000&&PE28_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE28.vbl=%b,value=%d@clk %d\n",PE28_Outport0[35:33],PE28_Outport0[31:0],i);
            end
            if(PE110_Outport0[35:33]!=3'b000&&PE110_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE110.vbl=%b,value=%d@clk %d\n",PE110_Outport0[35:33],PE110_Outport0[31:0],i);
            end
            if(PE6_Outport0[35:33]!=3'b000&&PE6_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE6.vbl=%b,value=%d@clk %d\n",PE6_Outport0[35:33],PE6_Outport0[31:0],i);
            end
            if(PE7_Outport0[35:33]!=3'b000&&PE7_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE7.vbl=%b,value=%d@clk %d\n",PE7_Outport0[35:33],PE7_Outport0[31:0],i);
            end
            if(PE8_Outport0[35:33]!=3'b000&&PE8_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE8.vbl=%b,value=%d@clk %d\n",PE8_Outport0[35:33],PE8_Outport0[31:0],i);
            end
            if(PE9_Outport0[35:33]!=3'b000&&PE9_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE9.vbl=%b,value=%d@clk %d\n",PE9_Outport0[35:33],PE9_Outport0[31:0],i);
            end
            if(PE29_Outport0[35:33]!=3'b000&&PE29_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE29.vbl=%b,value=%d@clk %d\n",PE29_Outport0[35:33],PE29_Outport0[31:0],i);
            end
            if(PE31_Outport0[35:33]!=3'b000&&PE31_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE31.vbl=%b,value=%d@clk %d\n",PE31_Outport0[35:33],PE31_Outport0[31:0],i);
            end
            if(PE10_Outport0[35:33]!=3'b000&&PE10_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE10.vbl=%b,value=%d@clk %d\n",PE10_Outport0[35:33],PE10_Outport0[31:0],i);
            end
            if(PE37_Outport0[35:33]!=3'b000&&PE37_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE37.vbl=%b,value=%d@clk %d\n",PE37_Outport0[35:33],PE37_Outport0[31:0],i);
            end
            if(PE11_Outport0[35:33]!=3'b000&&PE11_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE11.vbl=%b,value=%d@clk %d\n",PE11_Outport0[35:33],PE11_Outport0[31:0],i);
            end
            if(PE12_Outport0[35:33]!=3'b000&&PE12_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE12.vbl=%b,value=%d@clk %d\n",PE12_Outport0[35:33],PE12_Outport0[31:0],i);
            end
            if(PE13_Outport0[35:33]!=3'b000&&PE13_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE13.vbl=%b,value=%d@clk %d\n",PE13_Outport0[35:33],PE13_Outport0[31:0],i);
            end
            if(PE109_Outport0[35:33]!=3'b000&&PE109_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE109.vbl=%b,value=%d@clk %d\n",PE109_Outport0[35:33],PE109_Outport0[31:0],i);
            end
            if(PE100_Outport0[35:33]!=3'b000&&PE100_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE100.vbl=%b,value=%d@clk %d\n",PE100_Outport0[35:33],PE100_Outport0[31:0],i);
            end
            if(PE102_Outport0[35:33]!=3'b000&&PE102_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE102.vbl=%b,value=%d@clk %d\n",PE102_Outport0[35:33],PE102_Outport0[31:0],i);
            end
            if(PE103_Outport0[35:33]!=3'b000&&PE103_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE103.vbl=%b,value=%d@clk %d\n",PE103_Outport0[35:33],PE103_Outport0[31:0],i);
            end
            if(PE104_Outport0[35:33]!=3'b000&&PE104_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE104.vbl=%b,value=%d@clk %d\n",PE104_Outport0[35:33],PE104_Outport0[31:0],i);
            end
            if(PE14_Outport0[35:33]!=3'b000&&PE14_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE14.vbl=%b,value=%d@clk %d\n",PE14_Outport0[35:33],PE14_Outport0[31:0],i);
            end
            if(PE21_Outport0[35:33]!=3'b000&&PE21_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE21.vbl=%b,value=%d@clk %d\n",PE21_Outport0[35:33],PE21_Outport0[31:0],i);
            end
            if(PE15_Outport0[35:33]!=3'b000&&PE15_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE15.vbl=%b,value=%d@clk %d\n",PE15_Outport0[35:33],PE15_Outport0[31:0],i);
            end
            if(PE16_Outport0[35:33]!=3'b000&&PE16_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE16.vbl=%b,value=%d@clk %d\n",PE16_Outport0[35:33],PE16_Outport0[31:0],i);
            end
            if(PE17_Outport0[35:33]!=3'b000&&PE17_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE17.vbl=%b,value=%d@clk %d\n",PE17_Outport0[35:33],PE17_Outport0[31:0],i);
            end
            if(PE101_Outport0[35:33]!=3'b000&&PE101_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE101.vbl=%b,value=%d@clk %d\n",PE101_Outport0[35:33],PE101_Outport0[31:0],i);
            end
            if(PE19_Outport0[35:33]!=3'b000&&PE19_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE19.vbl=%b,value=%d@clk %d\n",PE19_Outport0[35:33],PE19_Outport0[31:0],i);
            end
            if(PE22_Outport0[35:33]!=3'b000&&PE22_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE22.vbl=%b,value=%d@clk %d\n",PE22_Outport0[35:33],PE22_Outport0[31:0],i);
            end
            if(PE23_Outport0[35:33]!=3'b000&&PE23_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE23.vbl=%b,value=%d@clk %d\n",PE23_Outport0[35:33],PE23_Outport0[31:0],i);
            end
            if(PE24_Outport0[35:33]!=3'b000&&PE24_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE24.vbl=%b,value=%d@clk %d\n",PE24_Outport0[35:33],PE24_Outport0[31:0],i);
            end
            if(PE111_Outport0[35:33]!=3'b000&&PE111_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE111.vbl=%b,value=%d@clk %d\n",PE111_Outport0[35:33],PE111_Outport0[31:0],i);
            end
            if(PE26_Outport0[35:33]!=3'b000&&PE26_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE26.vbl=%b,value=%d@clk %d\n",PE26_Outport0[35:33],PE26_Outport0[31:0],i);
            end
            if(PE27_Outport0[35:33]!=3'b000&&PE27_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE27.vbl=%b,value=%d@clk %d\n",PE27_Outport0[35:33],PE27_Outport0[31:0],i);
            end
            if(PE25_Outport0[35:33]!=3'b000&&PE25_Outport0[32]!=1'b1) begin
                $fwrite(filez,"PE25.vbl=%b,value=%d@clk %d\n",PE25_Outport0[35:33],PE25_Outport0[31:0],i);
            end
        end
        #1 $fclose(filez);
        $finish;
    end


  always #(CYCLE/2) clk=~clk;
endmodule
